 module Vote_test;
 wire[11:0] out;
 reg clk,Power,Close,Clear,Ballot,Total,Result;
 reg [3:0] IN;
 Vote v(clk,Power,Close,Clear,Ballot,Total,Result,IN,out);
 always #5 clk=~clk;
 initial begin
     Clear=1'b0;IN=3'b000;Close=1'b0;Total=1'b0;Result=1'b0;clk=1'b0;Ballot=1'b0;     
     #101 Power=1'b1;   
        #100 Clear=1'b1;#20 Clear=1'b0;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0010;#20 IN=4'b0000;
	#100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0101;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0101;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0101;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0101;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0101;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#200 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0011;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0011;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0011;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0010;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1000;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1000;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1111;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0010;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0011;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0011;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0011;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0011;#20 IN=4'b0000;#15 IN=4'b1000;#20 IN=4'b0000;#15 IN=4'b0011;#20 IN=4'b0000;
        #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1000;#20 IN=4'b0000;
	 #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1000;#20 IN=4'b0000;
	 #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1000;#20 IN=4'b0000;
	 #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1000;#20 IN=4'b0000;
	 #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1000;#20 IN=4'b0000;
	 #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1000;#20 IN=4'b0000;
	  #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1100;#20 IN=4'b0000;
	 #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1010;#20 IN=4'b0000;
	 #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1100;#20 IN=4'b0000;
	 #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1001;#20 IN=4'b0000;
	 #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1001;#20 IN=4'b0000;
	 #100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1001;#20 IN=4'b0000;
             
        #230 Total=1'b1;#34 Total=1'b0;
        #100 Close=1'b1;#22 Close=1'b0;
        
        #20 Result=1'b1; #20 Result=1'b0;
        #20 Result=1'b1; #20 Result=1'b0;
        #20 Result=1'b1; #20 Result=1'b0;
        #20 Result=1'b1; #20 Result=1'b0;
        #20 Result=1'b1; #20 Result=1'b0;
        #20 Result=1'b1; #20 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        
        #30 Clear=1'b1;#20 Clear=1'b0;
	#100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
	#100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0101;#20 IN=4'b0000;
	#100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b1111;#20 IN=4'b0000;
	#100 Ballot=1'b1;#25 Ballot=1'b0; #15 IN=4'b0001;#20 IN=4'b0000;
	#23 Total=1'b1;#34 Total=1'b0;
	#13 Close=1'b1;#32 Close=1'b0;
	#10 Power=1'b0;#20 Power=1'b1;
	#11 Close=1'b1;#22 Close=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
	#20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        #20 Result=1'b1; #45 Result=1'b0;
        #100 Clear=1'b1; Clear=1'b0;          
        #10 Power=1'b0;
        #100 Power=1'b1;
        #10 Ballot=1'b1;#30 Ballot=1'b0;
        #30 $finish;
 end
initial begin
    $dumpfile("V.vcd");
    $dumpvars(0,Vote_test);
    $monitor("Time=%d,Display=%d",$time,out);
end
 endmodule
